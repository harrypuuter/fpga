library verilog;
use verilog.vl_types.all;
entity teiler_vlg_vec_tst is
end teiler_vlg_vec_tst;
