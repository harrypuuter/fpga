library verilog;
use verilog.vl_types.all;
entity teiler is
    port(
        clock           : in     vl_logic;
        output          : out    vl_logic
    );
end teiler;
