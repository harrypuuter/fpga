library verilog;
use verilog.vl_types.all;
entity teiler is
    port(
        clock           : in     vl_logic;
        \out\           : out    vl_logic
    );
end teiler;
